module signExtend(i_data, o_data, enable);
input  [15:0]  i_data;
input [1:0] enable;
output reg [31:0]  o_data;

reg  [15:0]  data_r;
reg  [1:0] enable_r;
initial 
begin
enable_r = 1;

data_r = 0'b1111111111111111;
#150 enable_r = 0;
data_r = 0'b1111111111111111;
end
initial #300 $finish;


assign {i_data, enable} = {data_r, enable_r};

always @(enable,i_data)
begin
case (enable)
1: begin
 o_data[31:16] = {16{i_data[15]}};
 o_data[15:0] = i_data[15:0];
end

0:begin 
assign o_data[31:0] = i_data[15:0];
end
default: o_data[31:0] = i_data[15:0];
endcase

end
endmodule
